overkoepelend